module types

pub struct Object {

}