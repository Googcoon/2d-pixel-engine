module gui

pub fn temp(dir string) {
	println(dir)
}