module graphics

import gg
import gx

[params]
pub struct WindowOptions {

}

[heap]
struct Window {

}

fn InitWindow() &Window {
	
}