module graphics

import gg
import gx

struct Window {

}