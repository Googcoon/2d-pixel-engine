module vixel

pub struct Object {

}