module vixel

import gg.m4

